LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_arith.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY divide IS
    PORT (
        cl1 : IN STD_LOGIC;
        clk_divide : OUT STD_LOGIC
    );
END divide;

ARCHITECTURE fuc_d OF divide IS
BEGIN
    
END fuc_d;